module mynot(y,i);

input i;
output y;
wire y;

mynor G1 (y,i,i);

endmodule